module sbox (
    input   wire [5:0] in
    ,output wire [3:0] out
);

        always_comb// Valuta la combinazione con uno switch-case
          case (in)
            6'b000000: out = 4'b0010;
            6'b000001: out = 4'b1110;
            6'b000010: out = 4'b1100;
            6'b000011: out = 4'b1011;
            6'b000100: out = 4'b0100;
            6'b000101: out = 4'b0010;
            6'b000110: out = 4'b0001;
            6'b000111: out = 4'b1100;
            6'b001000: out = 4'b0111;
            6'b001001: out = 4'b0100;
            6'b001010: out = 4'b1010;
            6'b001011: out = 4'b0111;
            6'b001100: out = 4'b1011;
            6'b001101: out = 4'b1101;
            6'b001110: out = 4'b0110;
            6'b001111: out = 4'b0001;

            6'b010000: out = 4'b1000;
            6'b010001: out = 4'b0101;
            6'b010010: out = 4'b0101;
            6'b010011: out = 4'b0000;
            6'b010100: out = 4'b0011;
            6'b010101: out = 4'b1111;
            6'b010110: out = 4'b1111;
            6'b010111: out = 4'b1100;
            6'b011000: out = 4'b1101;
            6'b011001: out = 4'b0011;
            6'b011010: out = 4'b0000;
            6'b011011: out = 4'b1001;
            6'b011100: out = 4'b1110;
            6'b011101: out = 4'b1000;
            6'b011110: out = 4'b1001;
            6'b011111: out = 4'b0110;

            6'b100000: out = 4'b0100;
            6'b100001: out = 4'b1011;
            6'b100010: out = 4'b0010;
            6'b100011: out = 4'b1000;
            6'b100100: out = 4'b0001;
            6'b100101: out = 4'b1100;
            6'b100110: out = 4'b1011;
            6'b100111: out = 4'b0111;
            6'b101000: out = 4'b1100;
            6'b101001: out = 4'b0001;
            6'b101010: out = 4'b1101;
            6'b101011: out = 4'b1110;
            6'b101100: out = 4'b0111;
            6'b101101: out = 4'b0010;
            6'b101110: out = 4'b1000;
            6'b101111: out = 4'b1101;

            6'b110000: out = 4'b1111;
            6'b110001: out = 4'b0110;
            6'b110010: out = 4'b1001;
            6'b110011: out = 4'b1111;
            6'b110100: out = 4'b1100;
            6'b110101: out = 4'b0000;
            6'b110110: out = 4'b0101;
            6'b110111: out = 4'b1001;
            6'b111000: out = 4'b0110;
            6'b111001: out = 4'b1100;
            6'b111010: out = 4'b0011;
            6'b111011: out = 4'b0100;
            6'b111100: out = 4'b0000;
            6'b111101: out = 4'b0101;
            6'b111110: out = 4'b1110;
            6'b111111: out = 4'b0011;
        endcase
endmodule